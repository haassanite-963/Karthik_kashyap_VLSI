module full_adder()
{
    
}